module cross_bar_demux_buffer #(
) (
);

endmodule
