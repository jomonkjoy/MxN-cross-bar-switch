module cross_bar_switch #(
) (
);

endmodule
