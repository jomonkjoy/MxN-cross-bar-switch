module arbiter_mx1 #(
) (
);

endmodule
